module m2(
clk,out
);

input clk;
input in;
output out;
endmodule
